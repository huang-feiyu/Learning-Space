`ifndef and_n2t
  `include "and_n2t.sv"
`endif
`define xor_n2t 1

module xor_n2t(input a, input b, output out);

  assign out = a ^ b;

endmodule