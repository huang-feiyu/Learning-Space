`ifndef not_n2t
  `include "not_n2t.sv"
`endif
`define or_n2t 1

module or_n2t(input a, input b, output out);

  assign out = a | b;

endmodule
